library IEEE;
use IEEE.STD_LOGIC_1164.all;

-- To use the testbench in tb_pipo.vhd,
-- please make sure that your entity declaration
-- is consistent with line24~30 of tb_pipo.vhd.