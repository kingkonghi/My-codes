    Mac OS X            	   2   �      �    ��������                          ATTR       �   �   4                  �   $  com.apple.decmpfs       �     com.apple.lastuseddate#PS    fpmc  ��          2ݗ��Hu�k�5meԏ�a    gW�    